module pc(
	input addr,
	input clk,
	output addr_out
	);

	

endmodule // pc